library verilog;
use verilog.vl_types.all;
entity muxdecod_vlg_check_tst is
    port(
        Saida           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end muxdecod_vlg_check_tst;
