library verilog;
use verilog.vl_types.all;
entity Block3_vlg_check_tst is
    port(
        LEDR            : in     vl_logic_vector(0 downto 0);
        sampler_rx      : in     vl_logic
    );
end Block3_vlg_check_tst;
