library verilog;
use verilog.vl_types.all;
entity muxdecod_vlg_vec_tst is
end muxdecod_vlg_vec_tst;
