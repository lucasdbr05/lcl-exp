library verilog;
use verilog.vl_types.all;
entity Block8_vlg_vec_tst is
end Block8_vlg_vec_tst;
