library verilog;
use verilog.vl_types.all;
entity Block9_vlg_vec_tst is
end Block9_vlg_vec_tst;
