library verilog;
use verilog.vl_types.all;
entity Block12_vlg_vec_tst is
end Block12_vlg_vec_tst;
