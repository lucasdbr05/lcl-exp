library verilog;
use verilog.vl_types.all;
entity Block7_vlg_vec_tst is
end Block7_vlg_vec_tst;
