library verilog;
use verilog.vl_types.all;
entity Block5_vlg_check_tst is
    port(
        \OUT\           : in     vl_logic_vector(9 downto 0);
        sampler_rx      : in     vl_logic
    );
end Block5_vlg_check_tst;
