library verilog;
use verilog.vl_types.all;
entity Block1_vlg_check_tst is
    port(
        LEDR            : in     vl_logic_vector(1 downto 0);
        sampler_rx      : in     vl_logic
    );
end Block1_vlg_check_tst;
