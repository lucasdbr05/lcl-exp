library verilog;
use verilog.vl_types.all;
entity muxABC_vlg_vec_tst is
end muxABC_vlg_vec_tst;
